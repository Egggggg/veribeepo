module driver(
    i_clk,
    o_segments_drive,
    
);

endmodule